// Verilog Hello world 
module top(output wire D1);
assign D1 = 1'b0;

endmodule
