// Verilog Hello world 
module top(output wire D1, D2);
assign D1 = 1'b0;
assign D2 = 1'b1;

endmodule
